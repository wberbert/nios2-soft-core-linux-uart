// NIOS2_Design.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module NIOS2_Design (
		input  wire        clk_clk,                        //                        clk.clk
		input  wire        reset_reset_n,                  //                      reset.reset_n
		output wire [12:0] sdram_0_wire_addr,              //               sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                //                           .ba
		output wire        sdram_0_wire_cas_n,             //                           .cas_n
		output wire        sdram_0_wire_cke,               //                           .cke
		output wire        sdram_0_wire_cs_n,              //                           .cs_n
		inout  wire [31:0] sdram_0_wire_dq,                //                           .dq
		output wire [3:0]  sdram_0_wire_dqm,               //                           .dqm
		output wire        sdram_0_wire_ras_n,             //                           .ras_n
		output wire        sdram_0_wire_we_n,              //                           .we_n
		input  wire        uart_0_external_connection_rxd, // uart_0_external_connection.rxd
		output wire        uart_0_external_connection_txd  //                           .txd
	);

	wire  [31:0] nios2_data_master_readdata;                           // mm_interconnect_0:NIOS2_data_master_readdata -> NIOS2:d_readdata
	wire         nios2_data_master_waitrequest;                        // mm_interconnect_0:NIOS2_data_master_waitrequest -> NIOS2:d_waitrequest
	wire         nios2_data_master_debugaccess;                        // NIOS2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_data_master_debugaccess
	wire  [27:0] nios2_data_master_address;                            // NIOS2:d_address -> mm_interconnect_0:NIOS2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                         // NIOS2:d_byteenable -> mm_interconnect_0:NIOS2_data_master_byteenable
	wire         nios2_data_master_read;                               // NIOS2:d_read -> mm_interconnect_0:NIOS2_data_master_read
	wire         nios2_data_master_readdatavalid;                      // mm_interconnect_0:NIOS2_data_master_readdatavalid -> NIOS2:d_readdatavalid
	wire         nios2_data_master_write;                              // NIOS2:d_write -> mm_interconnect_0:NIOS2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                          // NIOS2:d_writedata -> mm_interconnect_0:NIOS2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                    // mm_interconnect_0:NIOS2_instruction_master_readdata -> NIOS2:i_readdata
	wire         nios2_instruction_master_waitrequest;                 // mm_interconnect_0:NIOS2_instruction_master_waitrequest -> NIOS2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                     // NIOS2:i_address -> mm_interconnect_0:NIOS2_instruction_master_address
	wire         nios2_instruction_master_read;                        // NIOS2:i_read -> mm_interconnect_0:NIOS2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;               // mm_interconnect_0:NIOS2_instruction_master_readdatavalid -> NIOS2:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;     // NIOS2:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;  // NIOS2:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;  // mm_interconnect_0:NIOS2_debug_mem_slave_debugaccess -> NIOS2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;      // mm_interconnect_0:NIOS2_debug_mem_slave_address -> NIOS2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;         // mm_interconnect_0:NIOS2_debug_mem_slave_read -> NIOS2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;   // mm_interconnect_0:NIOS2_debug_mem_slave_byteenable -> NIOS2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;        // mm_interconnect_0:NIOS2_debug_mem_slave_write -> NIOS2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;    // mm_interconnect_0:NIOS2_debug_mem_slave_writedata -> NIOS2:debug_mem_slave_writedata
	wire         mm_interconnect_0_mmu_s1_chipselect;                  // mm_interconnect_0:MMU_s1_chipselect -> MMU:chipselect
	wire  [31:0] mm_interconnect_0_mmu_s1_readdata;                    // MMU:readdata -> mm_interconnect_0:MMU_s1_readdata
	wire   [7:0] mm_interconnect_0_mmu_s1_address;                     // mm_interconnect_0:MMU_s1_address -> MMU:address
	wire   [3:0] mm_interconnect_0_mmu_s1_byteenable;                  // mm_interconnect_0:MMU_s1_byteenable -> MMU:byteenable
	wire         mm_interconnect_0_mmu_s1_write;                       // mm_interconnect_0:MMU_s1_write -> MMU:write
	wire  [31:0] mm_interconnect_0_mmu_s1_writedata;                   // mm_interconnect_0:MMU_s1_writedata -> MMU:writedata
	wire         mm_interconnect_0_mmu_s1_clken;                       // mm_interconnect_0:MMU_s1_clken -> MMU:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                  // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;               // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                   // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                      // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;             // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                     // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                 // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_timer_0_s1_chipselect;              // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                 // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                   // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;               // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                 // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                   // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                    // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                       // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;              // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                      // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                  // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;              // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                 // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                   // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;               // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_mmu_s2_chipselect;                  // mm_interconnect_0:MMU_s2_chipselect -> MMU:chipselect2
	wire  [31:0] mm_interconnect_0_mmu_s2_readdata;                    // MMU:readdata2 -> mm_interconnect_0:MMU_s2_readdata
	wire   [7:0] mm_interconnect_0_mmu_s2_address;                     // mm_interconnect_0:MMU_s2_address -> MMU:address2
	wire   [3:0] mm_interconnect_0_mmu_s2_byteenable;                  // mm_interconnect_0:MMU_s2_byteenable -> MMU:byteenable2
	wire         mm_interconnect_0_mmu_s2_write;                       // mm_interconnect_0:MMU_s2_write -> MMU:write2
	wire  [31:0] mm_interconnect_0_mmu_s2_writedata;                   // mm_interconnect_0:MMU_s2_writedata -> MMU:writedata2
	wire         mm_interconnect_0_mmu_s2_clken;                       // mm_interconnect_0:MMU_s2_clken -> MMU:clken2
	wire         irq_mapper_receiver0_irq;                             // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                             // uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                             // timer_1:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_irq_irq;                                        // irq_mapper:sender_irq -> NIOS2:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [JTAG:rst_n, MMU:reset, MMU:reset2, NIOS2:reset_n, SDRAM:reset_n, irq_mapper:reset, mm_interconnect_0:NIOS2_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, timer_0:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [MMU:reset_req, MMU:reset_req2, NIOS2:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                      // NIOS2:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                   // rst_controller_001:reset_out -> [mm_interconnect_0:timer_1_reset_reset_bridge_in_reset_reset, timer_1:reset_n]

	NIOS2_Design_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	NIOS2_Design_MMU mmu (
		.clk         (clk_clk),                             //   clk1.clk
		.address     (mm_interconnect_0_mmu_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_mmu_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_mmu_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_mmu_s1_write),      //       .write
		.readdata    (mm_interconnect_0_mmu_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_mmu_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_mmu_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),  //       .reset_req
		.address2    (mm_interconnect_0_mmu_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_mmu_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_mmu_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_mmu_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_mmu_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_mmu_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_mmu_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                             //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),      // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze      (1'b0)                                 // (terminated)
	);

	NIOS2_Design_NIOS2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	NIOS2_Design_SDRAM sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                        //  wire.export
		.zs_ba          (sdram_0_wire_ba),                          //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                       //      .export
		.zs_cke         (sdram_0_wire_cke),                         //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                        //      .export
		.zs_dq          (sdram_0_wire_dq),                          //      .export
		.zs_dqm         (sdram_0_wire_dqm),                         //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                       //      .export
		.zs_we_n        (sdram_0_wire_we_n)                         //      .export
	);

	NIOS2_Design_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	NIOS2_Design_timer_0 timer_1 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	NIOS2_Design_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_0_external_connection_rxd),          // external_connection.export
		.txd           (uart_0_external_connection_txd),          //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	NIOS2_Design_mm_interconnect_0 mm_interconnect_0 (
		.CLK_50_clk_clk                            (clk_clk),                                              //                          CLK_50_clk.clk
		.NIOS2_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                       //   NIOS2_reset_reset_bridge_in_reset.reset
		.timer_1_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   // timer_1_reset_reset_bridge_in_reset.reset
		.NIOS2_data_master_address                 (nios2_data_master_address),                            //                   NIOS2_data_master.address
		.NIOS2_data_master_waitrequest             (nios2_data_master_waitrequest),                        //                                    .waitrequest
		.NIOS2_data_master_byteenable              (nios2_data_master_byteenable),                         //                                    .byteenable
		.NIOS2_data_master_read                    (nios2_data_master_read),                               //                                    .read
		.NIOS2_data_master_readdata                (nios2_data_master_readdata),                           //                                    .readdata
		.NIOS2_data_master_readdatavalid           (nios2_data_master_readdatavalid),                      //                                    .readdatavalid
		.NIOS2_data_master_write                   (nios2_data_master_write),                              //                                    .write
		.NIOS2_data_master_writedata               (nios2_data_master_writedata),                          //                                    .writedata
		.NIOS2_data_master_debugaccess             (nios2_data_master_debugaccess),                        //                                    .debugaccess
		.NIOS2_instruction_master_address          (nios2_instruction_master_address),                     //            NIOS2_instruction_master.address
		.NIOS2_instruction_master_waitrequest      (nios2_instruction_master_waitrequest),                 //                                    .waitrequest
		.NIOS2_instruction_master_read             (nios2_instruction_master_read),                        //                                    .read
		.NIOS2_instruction_master_readdata         (nios2_instruction_master_readdata),                    //                                    .readdata
		.NIOS2_instruction_master_readdatavalid    (nios2_instruction_master_readdatavalid),               //                                    .readdatavalid
		.JTAG_avalon_jtag_slave_address            (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //              JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write              (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                    .write
		.JTAG_avalon_jtag_slave_read               (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                    .read
		.JTAG_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                    .readdata
		.JTAG_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                    .writedata
		.JTAG_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.JTAG_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.MMU_s1_address                            (mm_interconnect_0_mmu_s1_address),                     //                              MMU_s1.address
		.MMU_s1_write                              (mm_interconnect_0_mmu_s1_write),                       //                                    .write
		.MMU_s1_readdata                           (mm_interconnect_0_mmu_s1_readdata),                    //                                    .readdata
		.MMU_s1_writedata                          (mm_interconnect_0_mmu_s1_writedata),                   //                                    .writedata
		.MMU_s1_byteenable                         (mm_interconnect_0_mmu_s1_byteenable),                  //                                    .byteenable
		.MMU_s1_chipselect                         (mm_interconnect_0_mmu_s1_chipselect),                  //                                    .chipselect
		.MMU_s1_clken                              (mm_interconnect_0_mmu_s1_clken),                       //                                    .clken
		.MMU_s2_address                            (mm_interconnect_0_mmu_s2_address),                     //                              MMU_s2.address
		.MMU_s2_write                              (mm_interconnect_0_mmu_s2_write),                       //                                    .write
		.MMU_s2_readdata                           (mm_interconnect_0_mmu_s2_readdata),                    //                                    .readdata
		.MMU_s2_writedata                          (mm_interconnect_0_mmu_s2_writedata),                   //                                    .writedata
		.MMU_s2_byteenable                         (mm_interconnect_0_mmu_s2_byteenable),                  //                                    .byteenable
		.MMU_s2_chipselect                         (mm_interconnect_0_mmu_s2_chipselect),                  //                                    .chipselect
		.MMU_s2_clken                              (mm_interconnect_0_mmu_s2_clken),                       //                                    .clken
		.NIOS2_debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),      //               NIOS2_debug_mem_slave.address
		.NIOS2_debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),        //                                    .write
		.NIOS2_debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),         //                                    .read
		.NIOS2_debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),     //                                    .readdata
		.NIOS2_debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),    //                                    .writedata
		.NIOS2_debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),   //                                    .byteenable
		.NIOS2_debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),  //                                    .waitrequest
		.NIOS2_debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),  //                                    .debugaccess
		.SDRAM_s1_address                          (mm_interconnect_0_sdram_s1_address),                   //                            SDRAM_s1.address
		.SDRAM_s1_write                            (mm_interconnect_0_sdram_s1_write),                     //                                    .write
		.SDRAM_s1_read                             (mm_interconnect_0_sdram_s1_read),                      //                                    .read
		.SDRAM_s1_readdata                         (mm_interconnect_0_sdram_s1_readdata),                  //                                    .readdata
		.SDRAM_s1_writedata                        (mm_interconnect_0_sdram_s1_writedata),                 //                                    .writedata
		.SDRAM_s1_byteenable                       (mm_interconnect_0_sdram_s1_byteenable),                //                                    .byteenable
		.SDRAM_s1_readdatavalid                    (mm_interconnect_0_sdram_s1_readdatavalid),             //                                    .readdatavalid
		.SDRAM_s1_waitrequest                      (mm_interconnect_0_sdram_s1_waitrequest),               //                                    .waitrequest
		.SDRAM_s1_chipselect                       (mm_interconnect_0_sdram_s1_chipselect),                //                                    .chipselect
		.timer_0_s1_address                        (mm_interconnect_0_timer_0_s1_address),                 //                          timer_0_s1.address
		.timer_0_s1_write                          (mm_interconnect_0_timer_0_s1_write),                   //                                    .write
		.timer_0_s1_readdata                       (mm_interconnect_0_timer_0_s1_readdata),                //                                    .readdata
		.timer_0_s1_writedata                      (mm_interconnect_0_timer_0_s1_writedata),               //                                    .writedata
		.timer_0_s1_chipselect                     (mm_interconnect_0_timer_0_s1_chipselect),              //                                    .chipselect
		.timer_1_s1_address                        (mm_interconnect_0_timer_1_s1_address),                 //                          timer_1_s1.address
		.timer_1_s1_write                          (mm_interconnect_0_timer_1_s1_write),                   //                                    .write
		.timer_1_s1_readdata                       (mm_interconnect_0_timer_1_s1_readdata),                //                                    .readdata
		.timer_1_s1_writedata                      (mm_interconnect_0_timer_1_s1_writedata),               //                                    .writedata
		.timer_1_s1_chipselect                     (mm_interconnect_0_timer_1_s1_chipselect),              //                                    .chipselect
		.uart_s1_address                           (mm_interconnect_0_uart_s1_address),                    //                             uart_s1.address
		.uart_s1_write                             (mm_interconnect_0_uart_s1_write),                      //                                    .write
		.uart_s1_read                              (mm_interconnect_0_uart_s1_read),                       //                                    .read
		.uart_s1_readdata                          (mm_interconnect_0_uart_s1_readdata),                   //                                    .readdata
		.uart_s1_writedata                         (mm_interconnect_0_uart_s1_writedata),                  //                                    .writedata
		.uart_s1_begintransfer                     (mm_interconnect_0_uart_s1_begintransfer),              //                                    .begintransfer
		.uart_s1_chipselect                        (mm_interconnect_0_uart_s1_chipselect)                  //                                    .chipselect
	);

	NIOS2_Design_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
